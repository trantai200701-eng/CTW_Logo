VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO logo_from_pixels
  CLASS BLOCK ;
  FOREIGN logo_from_pixels ;
  ORIGIN -1.600 0.000 ;
  SIZE 48.000 BY 55.200 ;
  OBS
      LAYER met5 ;
        RECT 8.000 54.400 43.200 55.200 ;
        RECT 7.200 53.600 44.000 54.400 ;
        RECT 6.400 52.800 44.800 53.600 ;
        RECT 5.600 52.000 45.600 52.800 ;
        RECT 4.800 51.200 46.400 52.000 ;
        RECT 4.000 50.400 47.200 51.200 ;
        RECT 3.200 49.600 48.000 50.400 ;
        RECT 2.400 48.800 48.800 49.600 ;
        RECT 1.600 46.400 49.600 48.800 ;
        RECT 1.600 28.800 9.600 46.400 ;
        RECT 14.400 33.600 49.600 42.400 ;
        RECT 1.600 21.600 29.600 28.800 ;
        RECT 1.600 8.800 9.600 17.600 ;
        RECT 1.600 7.200 11.200 8.800 ;
        RECT 1.600 6.400 12.000 7.200 ;
        RECT 21.600 6.400 29.600 15.200 ;
        RECT 33.600 11.200 40.000 33.600 ;
        RECT 44.800 8.800 49.600 28.800 ;
        RECT 43.200 7.200 49.600 8.800 ;
        RECT 42.400 6.400 49.600 7.200 ;
        RECT 2.400 5.600 48.800 6.400 ;
        RECT 3.200 4.800 48.000 5.600 ;
        RECT 4.000 4.000 47.200 4.800 ;
        RECT 4.800 3.200 46.400 4.000 ;
        RECT 5.600 2.400 45.600 3.200 ;
        RECT 6.400 1.600 44.800 2.400 ;
        RECT 7.200 0.800 44.000 1.600 ;
        RECT 8.000 0.000 43.200 0.800 ;
  END
END logo_from_pixels
END LIBRARY

