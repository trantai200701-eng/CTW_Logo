magic
tech sky130A
timestamp 1762933526
<< metal5 >>
rect 800 5440 4320 5520
rect 720 5360 4400 5440
rect 640 5280 4480 5360
rect 560 5200 4560 5280
rect 480 5120 4640 5200
rect 400 5040 4720 5120
rect 320 4960 4800 5040
rect 240 4880 4880 4960
rect 160 4640 4960 4880
rect 160 2880 960 4640
rect 1440 3360 4960 4240
rect 160 2160 2960 2880
rect 160 880 960 1760
rect 160 720 1120 880
rect 160 640 1200 720
rect 2160 640 2960 1520
rect 3360 1120 4000 3360
rect 4480 880 4960 2880
rect 4320 720 4960 880
rect 4240 640 4960 720
rect 240 560 4880 640
rect 320 480 4800 560
rect 400 400 4720 480
rect 480 320 4640 400
rect 560 240 4560 320
rect 640 160 4480 240
rect 720 80 4400 160
rect 800 0 4320 80
<< end >>
